﻿"LOCATION","INDICATOR","SUBJECT","MEASURE","FREQUENCY","TIME","Value","Flag Codes"
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",2.496043,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",2.20621,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",2.06232,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",-1.605659,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",3.704804,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",1.664839,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",-0.11575,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",4.226493,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",0.513756,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.118313,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.884794,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",1.201876,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.740876,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.173227,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",-0.188855,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",0.05365,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.134519,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",-0.311348,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",0.329498,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.575565,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",2.28358,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.063471,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",0.216597,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",0.173414,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",2.997686,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.461092,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",3.387472,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",3.146134,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",0.863092,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",1.130646,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.501605,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.514168,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.300768,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",-0.329084,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.344931,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.505497,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.130099,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",3.444241,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.86505,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.655426,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.175864,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.410278,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.701658,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.441854,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",2.509552,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.271691,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.129321,
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.058315,"E"
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.23097,"E"
"AUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.077323,"E"
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-2.730124,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.175137,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.465527,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",1.368857,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.043233,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.876584,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-0.201445,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.201412,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",1.303772,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.781856,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.354356,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-5.043286,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.421345,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",1.784201,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.848736,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.020661,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.970912,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",2.497956,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.500765,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-3.380664,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-3.071392,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.18258,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",2.836727,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",2.660356,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.284889,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.779574,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.09776,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.726637,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.902228,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.250454,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.786519,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.423517,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.697084,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",2.400129,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.135251,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.862284,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.567644,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-3.478708,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",0.961438,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.754984,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.292667,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.548672,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.873736,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.216551,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-1.205697,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.984957,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.022829,
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.615358,"E"
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-2.711286,"E"
"AUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-0.901887,"E"
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.135982,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",0.873047,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",3.77043,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.765113,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.405277,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.268919,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.87146,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.83356,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.911383,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.451354,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.616501,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.563959,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.000638,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.706843,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.464726,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.021087,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.074056,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.662865,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.373354,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.417601,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.122908,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.212311,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.530617,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-0.122141,
"AUT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.172556,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",2.072648,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.095353,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-0.291606,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.562367,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.705186,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.38379,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.707594,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.33843,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.176546,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.879802,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.295884,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.802251,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.138482,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.311211,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.13188,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.548914,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.836004,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.230016,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.496085,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-1.385316,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.826363,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.398848,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.468707,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.158278,
"AUT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-9.119049,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",3.595608,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",6.960996,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",6.771718,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",4.281784,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",0.636895,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",6.052682,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",2.507903,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.749378,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.376932,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",5.851172,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.985559,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.795543,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",1.27213,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",1.061274,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",0.801257,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.375202,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.49359,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",3.468119,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.456162,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.165336,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",3.824619,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.125212,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.500034,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",3.666697,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",0.420792,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.247508,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.635866,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.713542,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.069466,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",0.794643,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.229044,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.68576,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.842988,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.231169,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.522921,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.518987,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.848551,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.614202,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.647906,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.518472,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-0.683018,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.497549,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.86254,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.432672,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.547212,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.097921,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",-0.196369,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.232198,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.724096,
"BEL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",3.1412,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.210431,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.959244,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.904195,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.38566,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.221738,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-0.539573,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.945667,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.955343,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-0.106176,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-1.396086,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-3.238979,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-2.220094,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.998418,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",1.380065,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.823314,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-0.5598,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.293628,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.865561,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.622967,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",1.662975,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-2.290669,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.948006,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-3.751085,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.719475,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.744523,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.12402,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.889665,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.021128,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.215243,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",2.648051,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.515589,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.564479,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.221855,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.103851,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.22899,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.355479,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.04792,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.275001,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.167374,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.395756,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.076622,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.382252,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.863977,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.30291,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.092638,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.658704,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.425671,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.121062,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.867933,
"BEL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-8.968611,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",2.46052,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",3.463108,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",2.383058,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",-0.005018,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",1.145191,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",5.895251,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",2.774885,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",0.736899,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",-0.984282,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",-0.294399,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",1.374247,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",1.380028,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.324938,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.717831,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",0.897458,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",-0.853768,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",0.462247,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",0.95846,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",0.239983,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",-0.112031,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",0.87922,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.045706,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.023288,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.987984,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.220932,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",-0.219905,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.807194,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.860241,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.526625,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.140329,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.595274,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.622386,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.248583,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",0.841961,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.220528,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.066713,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",-0.006323,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.284687,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",0.480315,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.017754,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.633932,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.218411,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.328163,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.622746,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.265081,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.163681,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.782451,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.319317,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.91764,
"CAN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",7.914436,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",0.171252,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",0.801109,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",3.081023,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",1.853636,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-1.140886,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.322678,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-0.525586,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",1.905564,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",3.710608,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",1.144371,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",0.820199,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-5.634418,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.716153,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",2.137426,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.861557,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",2.005531,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",2.237516,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",2.086584,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.256985,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-1.223483,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-4.138227,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-2.285973,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-0.47482,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",1.341572,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.410861,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.784097,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.416064,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.155735,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.740957,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.030008,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.8909,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.276972,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.637861,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.276918,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.013237,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.530206,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.09176,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.201669,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.486767,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.922902,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.499443,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.442623,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.073572,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.761742,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.176263,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.299035,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.028323,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.671484,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.504015,
"CAN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-12.879715,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.771364,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",6.193066,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.858222,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-0.280971,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.151408,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.987405,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.33184,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",7.677927,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.555754,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",5.176794,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",4.167527,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",5.193672,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",6.153752,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",4.239151,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.322283,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.313646,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.337742,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.678646,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.41426,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.319222,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.155667,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",5.229985,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.351676,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",3.425115,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.371441,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.699721,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.428349,
"CZE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",0.302391,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.08041,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.342252,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.542004,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.124641,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-0.423137,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-0.473954,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.217311,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-3.85228,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.243488,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.52316,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.568888,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.069403,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.258718,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.727207,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.961509,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.97411,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.150175,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.276537,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.31291,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.377548,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.958706,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.021974,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",2.681559,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.453083,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.44895,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.082233,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-6.46988,
"CZE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",3.048569,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",5.076012,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",5.310813,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",5.454614,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",0.641074,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",4.10963,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",3.694287,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.706802,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",2.867729,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",3.442676,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",-0.771006,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.943594,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.790723,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.979318,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.02289,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",2.529066,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.16796,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.030952,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.962466,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.093386,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.926287,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",2.613889,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",1.721754,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.910343,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",6.384333,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.488079,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.384178,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",0.724837,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",-0.115174,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.018541,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.316299,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",-0.353033,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.822161,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.650364,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.193264,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.368854,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.317917,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.184416,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-1.488722,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.921726,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.913554,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.346245,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.911281,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.786338,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.584132,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.427971,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.19061,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.869077,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.201011,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.441278,
"DNK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.766192,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-2.464769,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.885071,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-1.880894,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-2.200143,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-5.627145,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",1.88909,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-2.079704,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.935003,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.157191,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.172821,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-3.468823,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",0.948417,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.294233,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",1.169052,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.398632,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",2.537777,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-1.875475,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-1.99538,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-1.456922,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-1.563236,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-1.457575,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.098246,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-2.204467,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-1.312063,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.051083,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.107291,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",2.071652,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.988664,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.565284,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.075253,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.82149,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.705089,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.496363,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.74818,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.656643,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.22179,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.299196,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.384744,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.54323,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.389798,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.570113,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-2.022579,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.246663,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.497105,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.209176,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.194113,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.304882,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.706402,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.265801,
"DNK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-3.023538,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.908178,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",7.611696,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",5.919263,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",3.170209,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",6.235548,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",1.439594,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",2.497404,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.596796,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",6.204744,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",3.531527,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.02786,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.888871,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",4.038921,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.141274,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.417666,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",4.131733,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.123108,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",4.625767,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",3.899095,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.399086,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",0.777131,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.620165,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",5.455784,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",4.429437,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.765807,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.065657,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",3.087258,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",4.01618,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.27188,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.325613,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.906201,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.957666,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.076265,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.382789,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.923572,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.424257,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",3.213598,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-1.169248,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-4.429144,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.483048,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.385086,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-1.607245,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.368264,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.197484,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.813473,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.349147,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",2.516491,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-1.143051,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-0.151493,
"FIN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.105341,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-2.558826,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.489109,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.442249,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.468992,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-4.585525,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.379002,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-2.475288,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.937875,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.605337,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",1.478948,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",0.855078,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-0.345418,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.476422,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.439607,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-0.289774,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-1.642522,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.135704,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.272477,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.778774,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-2.122058,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-7.120579,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-7.197072,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-6.254942,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.87508,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",2.017566,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.236136,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",2.844265,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.115841,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.823777,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.178138,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.461634,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.498296,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.308704,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.296921,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.496046,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.175633,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.588695,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.502301,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.273651,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.742578,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.679285,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.262582,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.719128,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.989075,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.595195,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.181162,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.423586,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.16304,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.275188,
"FIN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-2.56265,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.971212,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",6.724341,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",5.773919,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",5.099046,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",1.200261,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",2.055696,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",4.690106,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",5.139402,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",3.053702,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.643325,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.335971,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",6.485311,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.432612,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.437981,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",4.019108,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.207972,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",0.98612,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",3.229434,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",3.564247,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.398493,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",1.25295,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.406914,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",0.930567,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.0634,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",2.486617,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.089627,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.654637,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.473556,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.441044,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.648651,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.871008,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.919445,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.570758,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.10513,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.887587,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.48965,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",-0.468669,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.638008,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.022803,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.294486,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.001301,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.326726,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.354258,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.9622,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.811302,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.279427,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",2.109769,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.409723,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.390128,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.353619,
"FRA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",-0.801698,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.617919,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-2.939765,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.263553,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-1.404593,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.588178,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",1.844931,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.61783,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.53674,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.043932,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.578102,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.795314,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-4.315393,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.69544,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-1.383857,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-2.789951,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-0.383325,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.010584,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.883213,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.154575,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.035533,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-0.699968,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.27926,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-1.971366,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.082994,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.730527,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.036113,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.312915,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.716934,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.428001,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.550581,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.615529,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-2.445711,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.456191,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.959546,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.014256,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.732372,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.273538,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.337451,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.371723,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.152723,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.685538,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.50243,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.278804,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.490006,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.106045,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.436642,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-0.247495,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.032426,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.100659,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-8.435858,
"FRA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",7.526755,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.364272,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.983052,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",5.100988,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",4.037166,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",3.762491,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",4.662283,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",4.118106,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.087135,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.863318,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",0.841889,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",1.662488,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",1.034649,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",3.281032,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.641189,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",2.307415,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",1.515231,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.367928,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",2.579541,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",3.480071,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",3.533561,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",3.476712,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.552646,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.947004,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.58796,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.506245,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.683218,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.450864,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.018347,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.135401,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.478991,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.51138,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.92708,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.769179,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",0.91072,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.578152,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.599242,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.18148,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.026011,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-3.01009,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.305172,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.600992,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.616968,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.474731,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.036425,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.509462,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.355337,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.782613,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.039718,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.36753,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.383302,
"DEU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",0.92735,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-1.982285,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.117299,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.612094,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-3.053214,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-4.097086,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.737684,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-0.547377,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",0.02993,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",1.222699,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.306637,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.259731,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.310395,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.386203,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",0.532256,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.249284,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.732051,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.002278,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.585524,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-0.314713,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",0.782668,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",0.803217,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.264539,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-3.403196,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.438347,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.160747,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-1.055144,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.696579,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.064903,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.773114,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.379876,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.882589,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.188661,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.423038,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.376454,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.688209,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.388746,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.001459,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.218565,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.427555,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",2.084881,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.301987,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.384633,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.309661,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.740117,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.107239,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.052134,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.505987,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.74241,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.458867,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.011741,
"DEU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",1.904306,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",5.768865,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",-0.848634,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",0.722781,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",-0.12829,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",3.153603,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",1.346772,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",-0.244348,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",3.429027,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",-2.000449,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",-3.361532,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.764991,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",2.048805,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.503301,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",5.001257,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",-0.527211,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",3.245046,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.424711,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",4.068949,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.849826,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",4.402424,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.054964,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",-2.837255,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.281291,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.614028,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-1.395971,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.587822,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-0.90761,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-7.049243,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-5.180475,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-2.28924,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-0.587963,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",3.576222,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-4.15505,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.403712,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-3.675869,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.28433,
"GRC","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.352639,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-4.030412,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.991007,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-0.53338,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-2.466148,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.73718,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.88279,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.45623,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-1.154857,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",2.008903,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",1.264422,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.221737,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.216273,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-1.056541,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.982355,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",3.868269,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-0.548663,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.068682,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.458873,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",1.662341,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",1.091516,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.694719,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",3.233418,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.011091,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.38689,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.807895,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.016345,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-4.736047,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-3.192525,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.47846,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.493985,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",1.746125,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-3.006222,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",4.260213,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-0.109923,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",5.762689,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.329513,
"GRC","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-11.014474,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",8.236426,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",6.075188,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",-1.852686,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",15.558086,"B"
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.380854,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.673392,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",3.457947,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",0.691327,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.910934,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",5.766682,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",5.688886,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.620115,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",6.000996,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",6.459919,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.252974,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.483487,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",2.644511,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-3.013026,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.295548,"B"
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.636219,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-1.288122,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.784427,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-1.173309,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.596625,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-2.268813,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",3.051503,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",4.050119,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.861208,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.994506,
"HUN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",-0.372639,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.494565,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-4.558087,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.239123,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-3.509668,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-1.160885,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.09853,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.993441,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-0.704774,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-1.375218,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-3.112382,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-6.755749,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-10.249822,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-5.997202,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",5.227779,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-12.752345,"B"
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.125903,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.650124,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.661224,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",2.653728,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.152498,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-1.374338,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.613998,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.736313,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.724312,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-1.838262,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.137372,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-2.001339,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.42339,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.544439,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.016082,"B"
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.474514,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.548701,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",1.292527,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",5.745583,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",2.316604,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",4.873366,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.450374,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.386874,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.712665,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-7.247921,
"HUN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",7.968256,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",10.079836,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.972352,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",4.931442,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",3.636868,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",0.139456,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",4.106445,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",11.00645,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",5.181505,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",4.937546,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",3.1567,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",-0.531436,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-0.541078,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",-3.041241,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.820571,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",-0.280055,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",3.477419,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.705465,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",2.501828,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.009763,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.734169,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",-0.377903,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",-3.373894,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",0.630998,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",4.520087,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",-1.948747,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.2869,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",4.201283,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",4.25618,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.590596,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",-0.190268,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.65334,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",4.171415,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.933946,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",7.820992,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",3.277476,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.804619,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",5.172177,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.061923,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",6.397169,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-1.027395,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.086141,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.144015,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.100473,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-0.044785,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.680352,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.109382,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.814014,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.560336,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.665756,
"ISL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.387594,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",1.717794,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.39052,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.305905,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",0.594681,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-0.741855,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.807962,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-2.714487,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.001154,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-1.03034,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",1.428224,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",3.622172,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",1.308339,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.377957,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",0.2337,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.76552,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.936643,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",4.503698,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-4.05853,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-2.829352,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-2.312397,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-1.078507,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.201825,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-0.344705,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-1.700232,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.574081,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.674741,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.757527,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.889057,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.149994,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",3.688943,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.92207,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-4.306385,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-2.300955,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-1.144869,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.610631,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.5496,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.770056,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-0.288797,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-13.16118,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.453645,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.439133,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.383341,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",1.421171,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.61415,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.655089,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",3.695358,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.945864,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.423121,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-3.352185,
"ISL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-8.364208,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",3.045228,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",8.761517,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",3.81687,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",4.47817,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",6.956357,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",2.561435,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",6.287128,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",6.961385,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",-0.951022,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",5.957134,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",5.186016,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",3.054365,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",1.136399,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",7.240634,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.185185,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",-1.465696,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",5.077533,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",4.757168,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",5.566767,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",4.495599,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",4.017572,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",5.01211,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.525791,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.424907,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",4.928802,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.997702,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",6.807088,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.089529,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",4.40956,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",5.202368,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.614082,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",5.310665,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.069942,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.916942,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.360871,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.576506,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.646137,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-2.784901,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",4.797473,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",11.667177,"B"
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.370897,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.420187,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-1.949857,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",5.038633,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",19.880842,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-1.187031,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",5.04818,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",5.264621,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.584677,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",9.228331,
"IRL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",7.267668,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.531996,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-3.578096,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.737126,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-1.837716,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.863147,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-2.699446,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",0.441265,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.059342,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",2.394231,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-3.659956,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-2.967343,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.803315,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-2.068716,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-3.353163,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-0.435057,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.024265,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.422528,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.780685,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.833811,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",3.918517,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-2.563117,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-2.391973,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-0.369774,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",2.906544,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",4.040685,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",2.539637,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",2.856047,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",5.100894,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",4.710741,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",2.636413,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",1.03994,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.183918,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.723926,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.983897,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",3.009077,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.69364,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.530881,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-3.845116,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-10.304808,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-9.288619,"B"
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-1.676951,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.879685,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",2.775466,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.77767,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",3.454164,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",2.110665,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.554231,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.333259,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.892743,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-4.111783,
"IRL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",4.982793,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.470421,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.953997,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",6.507835,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",5.537087,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-1.369485,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",6.168858,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",4.150103,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.45388,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",5.1631,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.899018,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.585723,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-0.401443,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",0.883193,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.806123,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",2.025823,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",1.695659,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.913289,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",2.888172,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",3.556383,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",0.963183,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",0.046264,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",1.399459,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.891467,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",4.200471,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",2.964617,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.114258,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.845539,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.068617,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",0.703256,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.871761,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.670605,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",-0.784174,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",-0.70863,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",0.838599,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.446789,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",-0.220154,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",-0.076009,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.570202,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.992054,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.273472,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.675089,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.534536,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.794849,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.079548,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.059368,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.307394,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.645094,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.012384,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.513879,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.256811,
"ITA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",-1.291065,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-2.992297,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.763061,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.099623,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.6871,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-1.321741,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.398783,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.943524,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.561492,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.466071,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",1.293468,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",0.121455,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",0.759118,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.246985,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.581141,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.72773,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.139359,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.24447,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",1.22054,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-0.237101,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",0.92842,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",1.390852,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.595202,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-2.752742,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-1.986837,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.077123,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.122749,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.06795,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.711662,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.899009,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.843933,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",1.205229,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.851627,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.309672,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.166026,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.214688,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.607867,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.948381,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.159465,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.914447,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.986469,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.313595,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-2.725928,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-2.809538,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.099102,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.870851,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.79915,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.206281,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.149199,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.234344,
"ITA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-10.599112,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.151312,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",8.385305,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",6.941608,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",2.162615,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",4.569062,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",2.35569,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.104367,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",4.549739,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",4.263001,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",2.351951,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",4.209142,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.540013,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.523539,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.414816,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",5.342485,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.572623,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",4.285659,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",5.639072,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",4.50105,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",5.100126,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",3.135856,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",1.450307,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.288781,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.342011,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",3.038309,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.595518,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.711473,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.120415,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.806259,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.892721,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.423018,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.84272,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.42531,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.288404,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.677295,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.160912,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.628057,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.290545,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.42147,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.091681,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.629424,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.094065,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.234727,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.177309,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",2.011117,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.100485,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.913891,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.553966,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.03935,
"JPN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.235358,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.462613,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.321063,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-1.285457,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-4.632641,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.61521,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.456039,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",0.260384,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.220455,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.332971,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.336315,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.665102,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",0.020679,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.396177,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",0.317808,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-0.786974,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.197579,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.127035,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.551752,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.031562,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.574259,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-0.020604,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.913931,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-2.975482,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.397108,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.6494,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.30483,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.954321,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-2.625444,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-3.236743,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.316615,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-1.256707,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.974817,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.075263,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.178209,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.108059,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.143781,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.738672,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-0.986752,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.325144,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.968963,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.436981,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.49699,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.053004,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.174542,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.322555,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.793039,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.935051,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.237997,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.050472,
"JPN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.328146,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",7.10319,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",2.948407,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",9.203657,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",5.129032,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",5.560662,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",6.859556,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",9.045154,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",6.202751,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",7.365386,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",-2.025796,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",4.064532,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",5.181033,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",11.696349,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",11.286854,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",4.843327,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",6.415117,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",8.022121,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",10.331033,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",6.738848,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",8.839943,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",8.224629,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",5.042123,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",4.944125,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",6.485155,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",6.276729,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",6.034919,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",6.604829,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",4.829684,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",9.241997,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.896175,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.360164,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",6.588994,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",4.640435,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",4.526781,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",4.704116,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.163364,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",6.327742,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",5.633284,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",3.458658,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",5.957468,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.893116,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.410712,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.245705,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.277111,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.365689,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.785021,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",4.466796,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",3.820278,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.363096,
"KOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",3.043604,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",1.198899,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",2.210412,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",3.369768,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",2.400397,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",0.453704,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",4.274755,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",1.425003,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",2.89874,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-0.307352,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-1.165618,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",1.463198,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",1.422174,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.018622,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-1.880078,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.848901,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",3.58037,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",3.3295,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.513854,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-0.674837,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.035734,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",1.349874,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",0.05644,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",0.812206,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",1.586517,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",2.109136,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.784626,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-1.337109,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-10.151375,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.314398,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",4.09786,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.668495,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.482578,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.935312,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.24179,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.588686,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.52912,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-0.999549,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-3.218096,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.076715,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.299316,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.002607,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.448994,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.440633,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.272433,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.891151,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.239494,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-1.528124,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-1.349851,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.313397,
"KOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-3.91436,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",-0.336012,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.973282,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",8.044938,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",2.746515,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-6.234009,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",1.702922,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.106834,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",5.748418,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.820194,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.104479,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.585604,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.477098,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",3.671231,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",6.469531,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",0.978295,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",7.990898,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.303027,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",4.010653,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",6.85829,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.06458,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",5.596744,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",0.384962,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.959834,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.442595,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",-1.823269,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.259182,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.601944,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.310608,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",3.482119,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",1.206498,"B"
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",-1.771475,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.764431,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.731034,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.856139,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.993978,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.078312,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.65428,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-4.828497,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.201848,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.684153,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-1.760898,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.391339,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.829405,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-0.248373,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.768374,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.989921,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",-1.480395,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-1.649991,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-0.029004,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.320091,
"LUX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",6.512587,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",2.050629,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",0.317404,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.867658,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",0.11288,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-1.442236,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.314521,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.681499,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.745556,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-0.708354,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.643908,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.400523,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.367251,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.685163,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.347172,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.629236,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.375465,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.949542,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",3.388454,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.744267,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",3.037169,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",1.503837,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",0.059223,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",0.759786,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.110219,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.87783,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.071938,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",2.426155,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",2.95466,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",3.046382,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",4.300242,"B"
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",3.772658,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",1.344155,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.610505,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.93756,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.091994,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.271548,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.600399,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",2.9326,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.793351,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.168062,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.50164,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.269168,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.250337,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.48319,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.057103,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.335241,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.625809,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.700328,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.203611,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.461905,
"LUX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",-1.206352,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",0.517426,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",-0.398271,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",-0.218903,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",-6.177797,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.130287,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-1.157159,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",5.88994,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-1.777079,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",5.884471,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.677585,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",-4.562878,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.12817,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.375601,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",-1.374607,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",3.249408,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.36903,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-3.299295,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.02023,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-4.976184,"B"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.805566,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.374984,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-0.478572,
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.546626,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.577446,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.393125,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.533542,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.471351,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-1.335775,"E"
"MEX","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-0.906902,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",1.377211,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",2.301788,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",3.527984,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-1.637746,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",4.052536,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",6.620901,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-1.976411,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",3.331516,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-2.058604,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-2.262316,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",3.426723,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-2.853814,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.318474,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",2.71773,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.041497,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-0.34396,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",3.185185,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-6.577464,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",9.21632,"B"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.38458,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",2.041354,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.683766,
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.812625,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.598717,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.164645,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.544492,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.670931,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.203712,"E"
"MEX","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-8.17818,"E"
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",5.127022,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",3.209913,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",6.630772,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",6.795347,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",3.361617,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",4.999276,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.086088,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",2.790437,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",1.246839,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.548877,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",-0.338088,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",1.170548,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",3.994104,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.763252,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",1.834406,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",1.364853,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.223512,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.812447,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.038552,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.446542,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",1.205998,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",-0.188535,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.603967,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.757237,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",-1.535089,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.369665,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.208025,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.455491,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.207117,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.232099,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.010131,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.729895,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.320404,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.724666,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.387927,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.487344,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.893447,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.574105,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.255694,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.065094,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.64084,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.148846,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.759906,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.740464,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.982921,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.155939,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.543902,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.32107,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-0.171196,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-1.139488,
"NLD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",2.208649,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-1.975942,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.69481,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-1.591175,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-3.134714,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-3.962947,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.020339,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.722189,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.039997,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.083425,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.856891,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.138812,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-2.826745,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-2.232789,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.092041,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.280407,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.853044,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",0.033073,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.938966,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.741317,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",2.003615,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",0.405538,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",1.133047,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-1.044819,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.58442,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",4.19067,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",2.64612,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.545575,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.531131,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",2.083465,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.210884,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.546056,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.143472,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.612607,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.095109,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.561267,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.782566,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.627873,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.19178,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-1.944587,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.215705,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.433064,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.249594,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.17239,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.313764,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.519727,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.810414,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.750742,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.088735,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.465068,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-3.230968,
"NLD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",1.983277,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",2.739141,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.80133,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",4.377859,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",1.041976,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-2.588116,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",-0.598538,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",-5.657893,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",1.362813,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",1.340251,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.970439,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",4.952775,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-0.337011,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",1.52176,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.374153,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",-1.508754,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",-2.633436,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",0.975607,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",5.788775,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",4.581304,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",3.527241,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",-1.765519,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.757666,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.390998,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",0.331987,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.037157,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.299455,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",3.315401,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",-1.5921,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.092927,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.013751,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.779539,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.944163,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.904212,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",-0.370668,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",-0.094404,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.375051,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",3.957445,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-3.284471,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",5.346065,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-0.872509,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.935429,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",3.750517,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-2.043003,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-0.074444,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",2.490877,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.980992,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.185494,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.263321,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-1.071782,
"NZL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.453064,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.533537,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.383996,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",1.26266,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",2.789939,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-0.918141,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.591566,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",1.434168,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.062327,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.551076,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.862453,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.694659,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",0.44419,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.582093,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",1.357356,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.72982,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-1.051936,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.173446,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-3.808541,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-4.430938,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-3.821281,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-3.637214,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-3.409938,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",2.795908,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",3.474042,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.920367,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.481168,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-1.486838,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.90558,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",3.491274,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-1.298565,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",1.122919,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",1.225186,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.701575,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",2.222892,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",2.276829,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.058076,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-1.040603,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.81083,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.171052,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.744789,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.024748,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.670162,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",3.186749,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",1.913278,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.218097,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",2.525014,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.153409,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.083154,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.279992,
"NZL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-3.524916,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",5.959463,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",6.050835,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",4.640242,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",3.745485,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",4.133877,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",5.539185,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.426482,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",4.359852,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",4.37246,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",2.052068,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.867829,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",0.894798,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",4.626726,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",5.597993,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.106533,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",1.017579,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.467933,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",0.087847,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",4.199811,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",3.366209,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",4.244126,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.130895,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.272651,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",3.730343,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",3.121607,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.24277,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.57257,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.077229,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.165781,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.820761,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.71467,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.22089,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.211398,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.025167,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.045614,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",-0.716818,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",-1.722569,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-2.964997,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",0.136359,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",0.425863,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-0.785877,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.856517,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.634939,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.722778,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.386871,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.577258,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.929739,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.488662,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-0.756749,
"NOR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.400044,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.960812,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.436714,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.808731,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.432173,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",0.232434,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-0.202026,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",0.286474,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.86229,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-0.343727,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",2.136064,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",0.380224,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.015732,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-0.937954,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",0.139219,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.05265,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",2.648172,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-0.197675,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-0.86379,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",-3.447008,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-1.712629,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-1.599448,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.132334,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-0.046397,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.693633,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.492824,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.218255,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",2.084763,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.943522,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.136748,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-1.235026,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-2.082615,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.282665,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-2.807958,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.306471,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.882414,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.29828,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.731284,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",2.265194,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.100537,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.955817,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.466147,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.491831,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.808934,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.114487,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.454719,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.391387,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-0.393856,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.945856,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.830664,
"NOR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-2.652276,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",4.94268,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",8.060385,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",4.09221,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",5.229877,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",4.692921,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",11.736274,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.584057,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",4.335674,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",5.496205,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",4.210127,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.806372,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.540623,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",3.138985,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.455804,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.602361,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",3.128084,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",6.743809,"B"
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",4.682568,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.209657,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.476828,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.343761,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.47065,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",4.042998,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",4.763241,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",6.134181,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",5.017332,
"POL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-1.711063,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.25232,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-1.084024,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.906363,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.150668,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-0.029163,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-6.303285,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.014471,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-2.936545,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-3.23205,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.586676,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.173048,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.987147,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.979346,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",4.539207,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",3.576067,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-1.237862,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.899337,"B"
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.048332,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.093078,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.263131,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.055552,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",3.826277,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.794016,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.077371,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.712111,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.189213,
"POL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-0.761308,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",5.401208,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",9.233479,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",12.750037,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",-4.933383,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-8.080223,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",6.09586,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",5.623946,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.677504,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",4.964643,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",2.881154,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",1.744587,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.802679,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",-4.047139,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",-1.034449,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.857707,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",4.595781,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.851728,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",4.797348,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.948523,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.366542,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",5.260021,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.582973,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",-0.132255,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",0.606587,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.449444,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.740289,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.967817,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.136772,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.208466,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",1.120463,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.0467,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.727053,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.437681,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.160593,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.130466,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.865629,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.557699,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.641138,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.408071,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.029783,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.529917,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.969223,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.406469,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-1.014138,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.01153,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.10612,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.794666,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.118854,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.470142,
"PRT","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.918733,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",2.056878,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.965904,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-1.408428,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",4.92116,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",0.181602,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-2.063419,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-1.077528,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.899543,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-0.430479,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.567451,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.97596,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.260532,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",3.588042,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-1.191835,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-1.228793,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-0.434841,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",3.60774,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",2.836073,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",3.714647,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",1.937179,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-0.565993,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-2.367957,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-2.022714,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.115183,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",2.501686,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.352684,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.929314,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",3.107708,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.088332,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.946479,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.178925,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.502769,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.731938,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.602536,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.528788,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.416331,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.736154,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-0.463342,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.817174,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.299922,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-3.035321,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-4.591485,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.759584,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.375022,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",2.226407,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",2.233094,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.941535,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",3.136926,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.170454,
"PRT","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-9.371123,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",6.361016,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",6.424159,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",5.036304,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.807747,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.218077,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.510397,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",7.18958,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",7.843855,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.830319,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",3.29951,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",5.983527,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",7.547393,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",2.155218,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.863061,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",6.443057,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.531141,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.531672,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.441522,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.987452,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",3.501032,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.367794,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",2.299265,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.339567,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.260667,
"SVK","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",4.921535,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.051423,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.64987,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-1.049556,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-2.91999,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-2.080068,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.144754,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-2.484655,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-2.186412,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",2.323474,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",3.127058,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",2.295405,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.946274,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",3.169881,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.882634,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.365344,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.686305,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.321064,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.86686,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.619289,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.585673,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.399932,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.525218,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.279644,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.203994,
"SVK","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-8.967717,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.098975,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",8.044277,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",6.317833,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",4.558431,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",1.702636,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",4.04505,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.700688,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",4.682848,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",4.064141,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",6.060233,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",4.17208,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",3.279381,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",3.917637,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",6.680654,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.964173,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",1.372381,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.180185,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.771968,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",1.857996,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",-0.131784,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",0.809883,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.823579,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.328305,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.928841,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",0.83637,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.107443,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-0.167184,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",-0.471206,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-0.352505,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",0.464861,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.16015,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.155111,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.297572,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",0.320567,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.390591,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.584805,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.105218,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.25753,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",2.409944,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.542173,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.476268,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.928561,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.442658,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.29786,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.791017,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.45087,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.871648,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.224332,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.167049,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-0.283257,
"ESP","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",-1.964619,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-0.394432,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.79606,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.47455,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",0.045573,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.165365,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.878351,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-2.003908,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-4.158952,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-4.720416,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-4.664227,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-4.718927,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-2.492837,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-2.52639,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-4.978197,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-1.941297,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.546239,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",4.059477,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",3.037801,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",2.715902,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",3.760528,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",1.542091,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-2.071314,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-3.494366,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.708151,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.757877,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.115123,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",3.446404,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",4.459284,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",4.455955,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",4.281847,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",3.227995,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.94391,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.796116,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.203277,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.348862,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.86918,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.488932,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.007068,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-6.806925,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.729114,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-2.620742,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-4.856888,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-2.47601,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",1.383346,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",3.120097,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",2.48113,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.901755,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.088882,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.10027,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-11.038589,
"ESP","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",7.106765,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",3.050682,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.401439,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",4.625577,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",2.36283,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",2.099313,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",-0.097122,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",0.309524,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",3.777377,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",3.251893,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",0.510472,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.878474,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",0.488353,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",1.013301,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.147013,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",0.901812,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.207247,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.879899,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",-0.106849,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",1.250457,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",0.043905,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",1.283052,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.212635,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.194914,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.51461,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.86511,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.716939,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",4.060313,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.642629,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.503721,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.633572,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.776103,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",3.571319,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.831817,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.478315,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.834767,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.924815,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.248504,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-1.741133,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.429882,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.505902,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.856622,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.512119,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.767296,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.171497,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",2.895448,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.598324,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.931869,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.328086,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.361114,
"SWE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.258393,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-2.708989,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-2.313145,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.811707,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",0.519602,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",0.064125,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.787256,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-2.244697,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-2.23646,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.339202,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.988641,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.539642,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",0.696102,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.82999,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",0.95253,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.089682,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.233542,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.108511,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",2.206268,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.706556,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.066139,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-3.055201,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-3.867215,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-4.726276,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.663647,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.498144,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.294431,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-1.00827,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.569971,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",2.622818,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.931258,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.397754,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.647624,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.831016,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.43392,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.376516,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.118564,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.420338,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.527735,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.775595,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",1.494503,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.548954,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.813454,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.429958,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.467596,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.48056,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.402855,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.260979,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.443063,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.371182,
"SWE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-3.895325,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",2.770808,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",3.011744,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",3.447918,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",3.07176,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-2.177585,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",1.720375,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.445387,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",0.193897,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.106168,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",3.063748,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",0.337027,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-1.193321,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",1.474761,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",3.122287,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",1.995897,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",0.08477,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",-0.784318,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",0.687825,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.491052,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.053344,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",-2.571488,"B"
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",0.885004,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",0.915702,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",0.700358,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.783982,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.164304,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.990062,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.230508,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-0.361003,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.250493,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.296452,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.583234,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",-0.489438,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",0.698293,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.436623,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.448426,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",2.008131,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.922451,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.023976,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.657529,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-0.467456,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.429224,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.876575,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.081218,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.64733,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.618826,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.826379,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.364134,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.623871,
"CHE","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.389965,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",0.051457,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.72566,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-0.999853,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-1.855886,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-4.383396,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.99671,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-0.713271,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.040713,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.0886,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",0.945894,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",0.568019,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-0.705451,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.049033,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.466216,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.206556,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.158872,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.675895,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",1.764545,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.015164,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",1.488402,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",0.460532,"B"
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.819713,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-1.680274,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-0.120455,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-2.156357,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-2.079592,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-0.989797,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.474832,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.576472,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.177685,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-1.19335,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.29076,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.28167,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.430287,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.156765,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.899348,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.043738,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.621557,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-1.175632,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.121158,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.434152,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.279887,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.196567,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.121945,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.161967,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.316102,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-1.163839,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.197874,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.131454,
"CHE","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-4.491213,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.246055,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.951683,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",1.805508,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",3.770506,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",6.7116,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",9.814435,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",1.042407,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",0.988562,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",-1.247735,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",-3.287561,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",4.353405,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.883099,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",4.370971,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",8.726142,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",1.087869,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",5.95492,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",9.351028,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.010171,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",-3.819745,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",7.499425,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",-3.106479,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.575516,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",12.316833,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",-10.959294,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",4.798439,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",3.126822,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",8.275499,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.115928,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-6.453037,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",8.518336,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",-5.960742,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",6.717922,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",6.599642,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",9.138561,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",6.317675,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.700407,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",5.313557,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.331874,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-4.124464,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.519722,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",5.498641,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.094364,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",6.751075,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-0.079091,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",4.091664,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.29842,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",4.757448,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.512585,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.911034,
"TUR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",6.81463,"E"
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-1.231891,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.170206,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",-1.073881,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.755491,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.178666,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.467152,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",0.248054,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-1.544579,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",-1.426355,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-1.190694,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.950663,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.81444,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.898001,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-4.264869,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.586159,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-1.302547,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",-1.579662,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-0.605265,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",2.455854,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.077711,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",2.424865,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",0.653885,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-5.345785,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",4.513519,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.710186,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",2.196047,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-2.158754,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.518505,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.941114,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-2.848247,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-1.155476,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.518104,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.961066,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.5942,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.263368,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.878966,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-1.48335,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-0.121995,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.088853,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",4.16727,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",3.867776,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",1.339082,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.32783,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",3.615799,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.564627,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.348817,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.297438,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.894144,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-4.285706,
"TUR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.621904,"E"
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",6.53356,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",5.901773,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",1.780976,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",-0.704842,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",-0.806779,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",4.432389,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",3.454957,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",4.775896,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",3.129457,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",1.007621,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",5.966412,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",2.960137,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",5.290786,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",-0.928588,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",1.149795,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.618105,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",3.693551,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",-0.158055,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",0.413896,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.075557,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",2.03267,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",4.766221,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",3.660132,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",2.449734,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.399683,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.477585,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",3.063671,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.369804,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.155156,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.466186,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.908632,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.586179,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.609263,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.242226,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.799434,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",2.101734,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.110825,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.039565,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.115195,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.486159,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.41463,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.672044,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.514658,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.088878,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",2.000321,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.265694,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.460652,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.451539,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.516394,
"GBR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.721189,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-3.357292,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-1.788817,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",4.42533,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-1.814896,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-0.654629,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",-1.43999,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",-0.918078,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",-0.524335,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.489855,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-3.163638,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-6.420381,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-0.819586,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-1.059159,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",3.057476,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",2.699554,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.288126,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.423948,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",5.691402,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.866635,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.618495,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-3.412503,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-4.409526,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-1.349971,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",1.103621,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.832312,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.695892,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.528666,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.488576,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.458285,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.144443,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.765103,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.875532,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.046348,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.571899,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.999589,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.211393,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.334377,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.015352,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.86483,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.138456,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.200431,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",1.482918,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.734233,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.117572,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.182632,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.695591,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.06658,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.590816,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.602957,
"GBR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-12.169775,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",3.750088,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",2.432212,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",2.373524,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",-0.902185,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",2.737749,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",2.422737,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",1.066948,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",0.79202,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",0.447863,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",0.020232,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.319752,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-0.321277,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.736349,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.084731,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",1.838955,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.262027,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",0.726712,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.15608,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",0.881018,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.712373,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",1.310106,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.43523,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",0.380736,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",0.847109,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",0.220025,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.486064,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.449522,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.249716,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.953948,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.746401,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.19397,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.766428,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.02378,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.616489,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",2.089042,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",0.946807,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.404249,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",1.280744,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",3.196011,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.642871,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.038302,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.377515,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.425423,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.375923,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.556997,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.302963,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.952882,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.054625,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.235405,
"USA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.57994,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-1.688008,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",1.666994,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",2.215199,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-0.554273,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-3.801583,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",1.902097,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",2.484404,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",3.605473,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",1.576014,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-1.424245,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-0.781227,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-2.423932,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.879562,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",4.130843,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",1.382836,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.258932,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.799232,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",2.054345,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",1.801004,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.948028,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-2.702484,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.237044,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",1.040652,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",1.91258,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",1.254665,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.08174,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.731244,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.999992,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.63113,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.193985,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-2.192138,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.979857,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.137917,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.294869,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.430392,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.856196,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-0.361781,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-2.068052,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-6.444915,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.754252,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.783542,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",1.181925,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.722858,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",1.177418,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.409592,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.649082,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.657005,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.306194,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.555285,
"USA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-6.297501,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",2.446232,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.007424,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",4.733136,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",1.350454,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",6.262574,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",7.242363,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",2.161109,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",5.968477,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",10.540309,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",7.005073,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",7.749171,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.214664,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.739191,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.155852,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.089662,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.886884,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.841234,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",4.684812,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",5.337028,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.120537,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",3.855318,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",2.203165,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",0.088357,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-3.370408,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.024546,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",4.56593,"B"
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.207551,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.613777,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.751703,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.44408,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",-0.057212,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.702617,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.960581,
"CHL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",13.571733,"E"
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",2.261373,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",4.446544,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",3.810352,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",0.644136,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-0.234569,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",2.832086,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",2.891682,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-1.960238,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-1.612092,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.997699,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-1.649708,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",2.708823,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-3.40636,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.192883,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.912061,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",1.071803,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",2.095153,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.326044,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.806073,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.22149,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-0.036734,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.299252,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.605064,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",8.475173,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",2.957139,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.334306,"B"
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.702881,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.953006,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.367405,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-1.01455,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-0.095605,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.349443,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.425479,
"CHL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-18.754352,"E"
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",5.802471,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",6.675845,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",5.065217,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",6.778739,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",5.918075,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",5.039397,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",7.547773,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-3.468884,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",2.096834,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",5.356103,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",-1.644894,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",3.329112,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.280434,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.575129,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.542858,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.625491,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",2.963227,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",5.818296,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.575365,
"EST","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",3.179068,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.808849,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.755121,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",3.030944,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.675213,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",3.969848,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",5.13385,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.610168,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.392452,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-16.213352,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.588776,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",9.352214,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.24158,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.55514,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.761105,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",2.603901,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.317909,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.770836,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-1.855421,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.071569,
"EST","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-6.235403,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",1.730838,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",0.544637,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",-0.812323,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",3.416442,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.717413,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",4.145567,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.875648,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",-1.274091,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",5.180995,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",2.491069,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",-0.570645,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",-0.660058,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",-1.361129,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",-1.014583,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.968092,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.097893,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.821282,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-0.104408,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",4.101714,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.914287,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",-1.829839,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.925895,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",4.586722,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.192185,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",3.677931,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.114107,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.134064,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.880407,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.91246,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",3.027723,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.306155,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.598992,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.056468,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.065559,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.730418,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.927298,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.613568,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.857944,
"ISR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",6.170373,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.138874,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",1.006741,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-0.033454,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",-1.158887,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",-0.311147,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.147647,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",-0.675309,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.158144,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.761302,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",1.211364,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",4.469012,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",1.115726,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",5.167287,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",4.098623,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",2.375186,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.216796,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-1.110235,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.017425,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.831744,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-3.15356,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.404214,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.614927,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-1.485722,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.088796,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.193644,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.041013,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.457739,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",0.255122,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.823581,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.563727,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.640179,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.236857,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.088235,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.330376,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.686826,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.447507,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.619329,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.997076,
"ISR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-9.480461,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",-2.14808,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.982457,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",-2.270326,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-2.124976,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",5.484289,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",5.112061,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.227332,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",7.067459,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",5.833756,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",5.191992,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",6.593516,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",5.843662,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",4.767544,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-4.509965,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.455973,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",2.750149,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.866662,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",2.077855,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.275221,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-2.692989,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.301006,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.676255,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.969791,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.143792,
"RUS","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",3.68077,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-3.311107,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",-7.52051,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-1.425299,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-1.348342,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-1.392036,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-2.985541,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",8.996678,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",4.763945,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.404992,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",2.934053,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",0.669095,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.676818,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.512236,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.796202,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.718412,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.502703,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.496351,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.967411,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.394404,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.955116,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.527925,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-1.316851,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.523189,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.289903,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.032607,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.149833,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.032534,
"RUS","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-6.201737,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",7.002656,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",7.780461,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.599866,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",3.627881,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.240788,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.490193,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.439374,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.0876,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.280005,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",6.75916,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",5.929375,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",4.293787,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.136131,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-6.310373,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.433142,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",3.629863,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-0.572536,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-0.978773,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.14416,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.557417,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",3.474614,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",3.762879,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.625993,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.601382,
"SVN","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.609922,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-3.607551,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-2.360382,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.864078,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.575366,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.131278,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.392381,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",2.893663,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.185865,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.994677,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-2.945826,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.522506,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",2.016016,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",3.491671,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-2.273024,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.362501,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-2.862061,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-2.265861,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.185873,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",1.4946,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.569708,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.33775,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.956341,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.44918,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.795254,
"SVN","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.433916,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.649088,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.467071,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.092669,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.256685,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.559348,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.611049,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.431588,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.015449,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",0.020546,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.549187,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.033221,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.414032,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",1.03208,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.79251,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.094855,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.546877,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.585053,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.011455,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.317996,
"OECD","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",3.181477,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.981383,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.589014,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.718823,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.378776,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.607121,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.86402,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.497179,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-0.364207,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.146828,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",0.874114,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.460273,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.350129,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.008405,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.712562,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.837881,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.697019,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.458352,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.759895,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-0.191221,
"OECD","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-7.818263,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.313377,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",2.308575,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.76915,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.16876,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.197654,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.067936,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.07644,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.333618,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.662892,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.129413,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.660825,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.959276,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.297872,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.302724,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.915813,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.545532,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.422189,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.901961,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.62368,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.430451,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.292359,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.586039,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.72852,
"EU28","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.730077,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",-1.523012,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",-0.454624,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.875658,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",-1.970623,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",-2.825339,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.882766,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",0.466554,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",1.074355,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",1.031597,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.700538,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",-1.183562,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.57577,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",0.059214,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",1.824051,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",0.535195,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",0.407157,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",1.032087,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",1.663083,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.815643,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",-0.459944,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-1.361671,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-1.404373,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",-1.147256,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",0.612412,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",0.383525,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.173373,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.643457,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",0.233894,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-0.049458,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.212258,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-1.22113,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.523,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.620324,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.290583,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.20444,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.918993,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",0.496653,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",-1.100472,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-4.776497,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.029953,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.432458,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",0.442849,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.015321,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.699278,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.607322,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.713067,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.588047,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.929009,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.21493,
"G-7","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-7.263358,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1971",4.13794,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1972",4.842423,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1973",4.19823,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1974",1.680805,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1975",2.129332,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",3.417048,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",2.767314,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",2.864779,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.220901,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",0.829678,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",2.621104,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",0.999638,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.736711,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.55022,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",2.703064,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.093117,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",1.8637,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",2.375967,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",2.270706,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.438588,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",1.79897,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",2.791261,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.550988,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.758387,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",1.460343,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.93157,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.892598,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.965903,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.584936,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.864478,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.850318,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",2.110539,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.872029,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.011333,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.713778,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.038965,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.930587,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.462083,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",0.557463,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.41025,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.729953,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.455742,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.930887,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.618405,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.953167,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.321926,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.199092,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.771168,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.059482,
"G-7","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",2.341545,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",4.026388,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",8.23277,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",8.323332,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",10.845565,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",8.225511,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",5.743204,"B"
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",7.511471,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-8.435719,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",2.693275,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",3.255903,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.153089,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",6.44345,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.070375,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.745935,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",4.410931,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.617985,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",4.225905,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.819241,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",4.464449,
"LVA","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.82345,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",3.520693,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.111651,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",1.066479,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-1.229784,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",3.408602,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",6.842703,"B"
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.081126,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",6.80194,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-15.10408,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-5.511367,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",4.320829,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",1.802746,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",2.994296,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.09993,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.348565,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.671176,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.052289,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.922163,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.225706,
"LVA","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-4.957366,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",4.322209,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",7.302979,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",5.493707,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",4.20211,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",1.243605,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",11.617329,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",4.710039,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",9.115209,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.413985,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",6.916062,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",7.997152,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",7.186417,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",2.377351,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-4.30976,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",4.081411,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",6.906079,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.040509,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",3.07927,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",1.892073,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",-0.769429,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-0.998277,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",7.384366,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.152294,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.913347,
"LTU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",5.909505,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.571278,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.684699,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",2.622266,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-4.452495,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",3.144711,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-3.772634,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",2.771261,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",2.155986,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",5.232699,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",2.418631,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.059792,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",4.89692,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.267751,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-10.009373,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.265269,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.454576,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",3.141393,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",1.47853,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.491867,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",3.787484,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",4.876803,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-1.521003,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.778264,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.902293,
"LTU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-5.730047,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.094209,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.866836,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.065054,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.381967,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",2.387501,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",1.490927,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.845745,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.485332,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.198285,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",0.887442,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.408893,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.902106,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.221512,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.102216,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.54496,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.501471,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.590134,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.930389,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.736858,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.083845,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.299033,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.513706,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.080299,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.591102,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",1.539079,
"EA19","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",0.044908,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.284681,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.532608,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.710529,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",1.301046,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",1.082603,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",0.333707,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-0.433945,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.380011,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.539897,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.230088,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.328867,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.522422,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.136442,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.739113,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.633096,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.068525,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.675151,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.311365,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.467739,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.648258,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.239766,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.85811,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.501271,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.692287,
"EA19","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-7.920678,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",4.350918,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",7.161331,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.512697,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",-3.065891,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",4.119881,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",4.693192,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-3.135748,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",2.74549,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",6.716335,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",0.367653,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.065197,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-0.008338,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.090676,
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",9.841706,"E"
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",-11.597074,"E"
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",-0.055432,"E"
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",-0.338194,"E"
"ZAF","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",0.420096,"E"
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-3.036635,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-5.046833,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",1.769577,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",7.280849,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.156389,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",-0.651813,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",4.959833,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-5.432163,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-4.721309,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",1.541501,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.208909,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",1.125932,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.392141,
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-9.110748,"E"
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",12.045058,"E"
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.142085,"E"
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.152008,"E"
"ZAF","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.516715,"E"
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",1.064395,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",1.824573,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",-1.064712,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",2.028292,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",0.398494,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-1.424604,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.106776,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.312018,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",1.802835,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",-0.588318,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",0.679352,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",1.409289,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.504043,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",-1.740078,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",3.944701,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.360772,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",3.150387,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",2.834583,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",11.682433,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",4.80069,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",-1.394062,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",5.231701,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.542483,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",3.215565,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",4.38458,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",2.358197,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.292773,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",2.511722,
"CRI","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",15.483893,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",0.418543,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",0.04165,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",2.069926,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",-5.917132,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",5.688775,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",2.905339,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",2.629401,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",-0.802175,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-1.552225,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",4.274238,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",3.473566,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-0.554159,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.152695,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",1.91229,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.922232,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",1.394205,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.25773,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",4.14646,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.644316,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",5.294745,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.106163,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-5.058319,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-7.248948,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-1.3119,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",4.973006,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-3.838155,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",-0.301541,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-0.803786,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-1.363798,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.588592,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.377044,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-1.406075,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-17.793426,
"CRI","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",12.778089,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",3.122068,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",-2.556818,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-3.685135,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-2.642533,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-3.614575,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",3.191403,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.75854,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",2.879407,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",4.609038,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",2.933926,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",3.604919,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.730512,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",5.276153,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.977397,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-3.314177,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",0.197528,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.883805,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.160073,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.883591,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",1.012979,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.153147,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.518366,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.699117,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",1.089299,
"BGR","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-4.142252,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",2.547758,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-11.323629,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",8.481724,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-5.380727,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",9.046628,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.878702,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",5.66779,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",2.884611,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",2.372372,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",4.559364,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",3.633773,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",3.284612,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",1.27865,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",1.242934,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",5.731131,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",4.478663,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",3.285923,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",-0.162236,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.653041,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",3.046257,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.582152,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",0.972677,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.710657,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.643515,
"BGR","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.34502,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",6.07918,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",6.106278,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",2.519559,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-0.926924,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.176408,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",3.746589,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",4.949225,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",3.025118,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",3.270687,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",3.367436,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.695063,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",1.683525,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.224591,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-6.525517,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",1.93804,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",4.166086,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.241059,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",3.317836,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",-1.994099,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",4.797496,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",2.845111,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.539265,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",1.000632,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",-1.054288,
"HRV","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-6.779292,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",1.282074,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.513411,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-0.244776,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.484133,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",4.713941,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.86762,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",0.73769,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",2.42465,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.786718,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.835049,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",3.157306,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.182041,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",2.169036,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-0.703937,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-2.903329,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-3.780492,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-4.107476,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-3.232089,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",2.123645,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-1.515204,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.526057,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",2.89667,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",2.851407,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",5.192963,
"HRV","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-0.97731,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",5.191562,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",-5.60333,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.091837,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",1.354932,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.094692,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",6.376413,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",16.738429,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",4.067816,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",11.99922,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",5.528814,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",8.143543,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",5.484849,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",11.100721,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-0.866794,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",-2.043293,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",3.840978,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",2.688541,"B"
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",4.984811,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",3.625081,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",4.669416,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",4.529363,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",6.176291,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",4.313345,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",3.992513,
"ROU","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",-2.182775,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-0.900091,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",1.074815,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-2.902171,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-1.512474,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",-0.513379,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.970426,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-6.392795,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-1.196927,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-0.839649,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",-0.200645,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",0.487415,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",3.170845,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.039264,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.893854,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-1.312144,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-1.380449,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-0.197572,"B"
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-0.8027,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.346883,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",-1.171778,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",0.754873,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",1.662129,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",0.752154,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.709802,
"ROU","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-1.360795,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.292042,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.942532,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",1.741632,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",2.122671,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",3.228112,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",2.052185,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",1.954651,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.933511,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",1.614116,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.122284,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",1.650795,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",0.937299,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",-0.261931,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-1.168566,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",2.977575,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",1.787611,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",0.53979,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",0.920276,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",0.673336,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",1.38326,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",0.456422,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.743675,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",0.702154,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",1.002917,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",0.598307,
"EU27_2020","GDPCAPCONTR","LPRDTY","AGRWTH","A","2021",0.220969,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",0.328446,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.577591,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",1.126855,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",0.674854,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",0.415195,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.060142,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",-1.068264,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",-0.439859,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",0.536541,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",0.370355,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",1.460803,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.81651,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",0.566633,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",-3.472757,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",-0.924762,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",-0.092503,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",-1.415449,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",-1.055796,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.759262,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.683492,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",1.314655,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",0.887062,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",1.174583,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",0.60672,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-6.581227,
"EU27_2020","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2021",5.161161,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1976",1.766699,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1977",0.008823,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1978",5.992244,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1979",2.875684,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1980",2.439707,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1981",-1.510308,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1982",-0.099158,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1983",2.087438,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1984",2.522221,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1985",0.798877,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1986",2.535289,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1987",0.868451,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1988",1.216528,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1989",-0.716092,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1990",2.070437,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1991",-3.537575,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1992",3.102524,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1993",-0.963362,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1994",1.019356,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1995",0.787553,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1996",1.010114,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1997",1.27581,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1998",0.734305,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","1999",-3.774826,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2000",-3.748455,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2001",0.391285,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2002",-2.146656,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2003",0.193679,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2004",5.806281,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2005",1.789345,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2006",6.434405,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2007",4.193745,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2008",0.115508,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2009",-2.611671,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2010",0.464188,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2011",3.437117,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2012",1.151275,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2013",3.642228,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2014",2.641478,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2015",0.945013,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2016",1.880426,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2017",1.692382,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2018",2.276295,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2019",4.578224,
"COL","GDPCAPCONTR","LPRDTY","AGRWTH","A","2020",21.116367,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1971",0.342035,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1972",0.470783,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1973",0.5547,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1974",0.574754,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1975",2.768873,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1976",0.527022,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1977",1.842412,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1978",0.066461,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1979",0.173087,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1980",-0.613208,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1981",1.702459,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1982",-1.04318,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1983",-2.583413,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1984",-1.714394,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1985",3.601454,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1986",1.061518,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1987",2.552043,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1988",1.147309,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1989",2.177823,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1990",0.219262,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1991",4.4156,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1992",-0.78223,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1993",4.73209,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1994",2.707409,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1995",2.778171,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1996",-1.002062,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1997",0.397488,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1998",-1.527758,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","1999",-2.826592,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2000",5.07014,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2001",-0.00377,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2002",3.436904,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2003",2.434702,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2004",-1.662522,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2005",1.624695,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2006",-0.923442,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2007",1.233891,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2008",1.954852,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2009",2.641069,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2010",2.805948,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2011",2.200164,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2012",1.552271,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2013",0.285705,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2014",0.662325,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2015",0.853521,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2016",-0.907611,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2017",-1.41926,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2018",-0.801649,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2019",-2.291076,
"COL","GDPCAPCONTR","LUTILISATION","AGRWTH","A","2020",-23.849597,
